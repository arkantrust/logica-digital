LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

----------------------------------------------------------

ENTITY CONTROLADOR IS

PORT(
  RX_DATA : IN STD_LOGIC_VECTOR(7 DOWNTO 0); --SALIDA A
  LEDS : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
);

END CONTROLADOR;

----------------------------------------------------------

ARCHITECTURE BEHAVIORAL OF CONTROLADOR IS
  SIGNAL WIRE1 : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
  PROCESS(RX_DATA, WIRE1)
  BEGIN
    CASE RX_DATA IS
      WHEN "00000011" => WIRE1 <= "0111"; --3
      WHEN "00000101" => WIRE1 <= "0011"; --5
      WHEN "00100111" => WIRE1 <= "0001"; --7
      WHEN "00001111" => WIRE1 <= "0000"; --15
      WHEN OTHERS => WIRE1 <= "1111";
    END CASE;
  END PROCESS;

  LEDS <= WIRE1;
END ARCHITECTURE BEHAVIORAL;